// Code your design here
`include "fifo.v"