// Code your testbench here
// or browse Examples
`include "tb.sv"